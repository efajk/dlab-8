//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:     
// Design Name: 
// Module Name:   BullandCow  
// Project Name:  
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module BullandCow(  
  input wire iCLK_50, reset,
	input PS2_CLK,
	input PS2_DATA,
	output wire oHS, oVS,
  output wire  oVGA_R,
  output wire  oVGA_G,
  output wire  oVGA_B,
	output wire [7:0] oLED
);









endmodule